`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:48:27 01/25/2025 
// Design Name: 
// Module Name:    fadder1bit_verilog 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fadder1bit_verilog(
    input a,
    input b,
    input cin,
    output sum,
    output cout
    );


endmodule
